module forwarding_unit (
    ADDR1, ADDR2, WB_ADDR, MEM_ADDR, EXE_ADDR, OP1SEL, OP2SEL, OPCODE,
    DATA1IDSEL, DATA2IDSEL, DATA1EXESEL, DATA2EXESEL, DATAMEMSEL
);

// Declaring input output ports
input [4:0] ADDR1, ADDR2, WB_ADDR, MEM_ADDR, EXE_ADDR;
input OP1SEL, OP2SEL;
input [6:0] OPCODE;
output DATA1IDSEL, DATA2IDSEL, DATAMEMSEL;
output [1:0] DATA1EXESEL, DATA2EXESEL;

// check OPCODE for store
wire STORE;
nand store(STORE, !OPCODE[6], OPCODE[5], !OPCODE[4], !OPCODE[3], !OPCODE[2], OPCODE[1], OPCODE[0]);


wire [4:0] WB_EXE_XNOR_DATA1, WB_EXE_XNOR_DATA2;
wire WB_EXE_DATA1, WB_EXE_DATA2;


assign WB_EXE_XNOR_DATA1 = (MEM_ADDR ~^ ADDR1);
assign WB_EXE_XNOR_DATA2 = (MEM_ADDR ~^ ADDR2);
assign WB_EXE_DATA1 = (WB_EXE_XNOR_DATA1[4] & WB_EXE_XNOR_DATA1[3] & WB_EXE_XNOR_DATA1[2] & WB_EXE_XNOR_DATA1[1] & WB_EXE_XNOR_DATA1[0]);
assign WB_EXE_DATA2 = (WB_EXE_XNOR_DATA2[4] & WB_EXE_XNOR_DATA2[3] & WB_EXE_XNOR_DATA2[2] & WB_EXE_XNOR_DATA2[1] & WB_EXE_XNOR_DATA2[0] & STORE);


wire [4:0] WB_ID_XNOR_DATA1, WB_ID_XNOR_DATA2;


assign WB_ID_XNOR_DATA1 = (WB_ADDR ~^ ADDR1);
assign WB_ID_XNOR_DATA2 = (WB_ADDR ~^ ADDR2);
assign DATA1IDSEL = (WB_ID_XNOR_DATA1[4] & WB_ID_XNOR_DATA1[3] & WB_ID_XNOR_DATA1[2] & WB_ID_XNOR_DATA1[1] & WB_ID_XNOR_DATA1[0]);
assign DATA2IDSEL = (WB_ID_XNOR_DATA2[4] & WB_ID_XNOR_DATA2[3] & WB_ID_XNOR_DATA2[2] & WB_ID_XNOR_DATA2[1] & WB_ID_XNOR_DATA2[0]);


wire [4:0] MEM_EXE_XNOR_DATA1, MEM_EXE_XNOR_DATA2;
wire MEM_EXE_DATA1, MEM_EXE_DATA2;

assign MEM_EXE_XNOR_DATA1 = (EXE_ADDR ~^ ADDR1);
assign MEM_EXE_XNOR_DATA2 = (EXE_ADDR ~^ ADDR2);
assign MEM_EXE_DATA1 = (MEM_EXE_XNOR_DATA1[4] & MEM_EXE_XNOR_DATA1[3] & MEM_EXE_XNOR_DATA1[2] & MEM_EXE_XNOR_DATA1[1] & MEM_EXE_XNOR_DATA1[0]);
assign MEM_EXE_DATA2_AND_INPUT = (MEM_EXE_XNOR_DATA2[4] & MEM_EXE_XNOR_DATA2[3] & MEM_EXE_XNOR_DATA2[2] & MEM_EXE_XNOR_DATA2[1] & MEM_EXE_XNOR_DATA2[0]);
assign MEM_EXE_DATA2 = (STORE & MEM_EXE_DATA2_AND_INPUT);

assign DATA1EXESEL[1] = (WB_EXE_DATA1 | MEM_EXE_DATA1);
assign DATA1EXESEL[0] = ((OP1SEL & WB_EXE_DATA1) | MEM_EXE_DATA1);

assign DATA2EXESEL[1] = (WB_EXE_DATA2 | MEM_EXE_DATA2);
assign DATA2EXESEL[0] = ((OP2SEL & WB_EXE_DATA2) | MEM_EXE_DATA2);

assign DATAMEMSEL = MEM_EXE_DATA2_AND_INPUT;

endmodule